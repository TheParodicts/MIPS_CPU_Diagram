module Encoder (
  input[31:0] Instruction,
  output [6:0] State_Sel
);
  reg[6:0] state_tmp;
  
  assign State_Sel = state_tmp; 
  
  always @(*)
    begin
      casez(Instruction)
        // 32'b000000xxxxxxxxxxxxxxxxxxxx100000: //ADD
        
        32'b000000????????????????????100001: //ADDU
          state_tmp = 7'd5;
        
        32'b101000??????????????????????????: //SB
          state_tmp = 7'd6;
        
        32'b000100??????????????????????????: //BEQ
          state_tmp = 7'd10;
        
        default: state_tmp = 7'd0;
      
      endcase      
    end
endmodule
